module uart_rx(
  input  wire        clock,
  input  wire        reset,
  input  wire        rx,
  output reg   [7:0] data,
  output reg         busy);
  
endmodule
